//----------------------------------------------------------------------
// CounterVRTL.v
//----------------------------------------------------------------------

`ifndef COUNTER_COUNTER_VRTL_V
`define COUNTER_COUNTER_VRTL_V


module CounterVRTL(
    input  logic        clk,
    input  logic        reset,
    input  logic        en,
    output logic [31:0] out
);

//----------------------------------------------------------------------
// SECTION TASK:
// Implement your design here
//----------------------------------------------------------------------



endmodule

`endif // COUNTER_COUNTER_VRTL_V